/*------------------------------------------------------------------------------
 * File          : oflow_define.txt
 * Project       : RTL
 * Author        : epchof
 * Creation date : Jan 6, 2024
 * Description   :
 *------------------------------------------------------------------------------*/



`define W_IOU_ADDR  3'h0 
`define W_WIDTH_ADDR  3'h1
`define W_HEIGHT_ADDR  3'h2
`define W_COLOR1_ADDR  3'h3
`define W_COLOR2_ADDR  3'h4
`define W_HISTORY_ADDR  3'h5
`define NUM_OF_HISTORY_FRAMES_ADDR 3'h6

`define ADDR_LEN 3