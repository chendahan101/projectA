/*------------------------------------------------------------------------------
 * File          : oflow_define.txt
 * Project       : RTL
 * Author        : epchof
 * Creation date : Jan 6, 2024
 * Description   :
 *------------------------------------------------------------------------------*/



`define W_IOU_ADDR  4'h0 
`define W_WIDTH_ADDR  4'h1
`define W_HEIGHT_ADDR  4'h2
`define W_COLOR1_ADDR  4'h3
`define W_COLOR2_ADDR  4'h4
`define W_HISTORY_ADDR  4'h5

`define SCORE_TH_FOR_NEW_BBOX_ADDR 4'h6
`define NUM_OF_HISTORY_FRAMES_ADDR 4'h7
`define MAX_THRESHOLD_FOR_CONFLICTS_ADDR 4'h8

`define ADDR_LEN 4