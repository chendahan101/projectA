/*------------------------------------------------------------------------------
 * File          : oflow_pe_conflict_resolve_fsm.sv
 * Project       : RTL
 * Author        : epchof
 * Creation date : Jun 27, 2024
 * Description   :
 *------------------------------------------------------------------------------*/

module oflow_pe_conflict_resolve_fsm #() ();

endmodule