/*------------------------------------------------------------------------------
 * File          : oflow_similarity_metric_define.sv
 * Project       : RTL
 * Author        : epchof
 * Creation date : Jun 13, 2024
 * Description   :
 *------------------------------------------------------------------------------*/


`include "/users/epchof/Project/design/work/include_files/oflow_MEM_buffer_define.sv"

`define BBOX_VECTOR_SIZE 89
`define MAX_BBOXES_PER_FRAME 256

`define REGISTER_DATA_LEN 10 // explenation in ipad, q0.9
`define REGISTER_ADD_LEN 10 // explenation in ipad, q0.9


`define ID_LEN 12

