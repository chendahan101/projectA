/*------------------------------------------------------------------------------
 * File          : oflow_MEM_buffer_define.sv
 * Project       : RTL
 * Author        : epchof
 * Creation date : Jun 23, 2024
 * Description   :
 *------------------------------------------------------------------------------*/
`define TOTAL_FRAME_NUM_WIDTH 8
`define NUM_OF_HISTORY_FRAMES_WIDTH 3
`define NUM_OF_BBOX_IN_FRAME_WIDTH 8
`define DATA_WIDTH 290
`define OFFSET_WIDTH 8
`define ADDR_WIDTH 8
